//Divider Stage Module and Pipelined Divider Module
