//testbench for pipelined divider
