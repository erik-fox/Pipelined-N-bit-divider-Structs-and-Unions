package mips;
  
  typedef union packed{
    struct packed {
    }r;
    struct packed {
    }i;
    struct packed {
    }i;
  }mipsinst;
endpackage
