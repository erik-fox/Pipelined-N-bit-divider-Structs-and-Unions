task sendByte();

endtask

task sendSegmentHeader();

endtask
